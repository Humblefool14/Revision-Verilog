always@(a,b)
  begin 
    sum = a+b;
    sub = a-b;
    prod = a*b;
  end 
