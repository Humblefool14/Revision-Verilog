  ahb_burst_e trans_burst[8] = '{AHB5_SINGLE,AHB5_INCR,AHB5_WRAP4, AHB5_INCR4, AHB5_WRAP8, AHB5_INCR8, AHB5_WRAP16, AHB5_INCR16};
