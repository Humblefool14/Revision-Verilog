

function new(string name = "AHBTXN");
    super.new(name);
  endfunction

  function void pre_randomize();
  endfunction

  function void post_randomize();
  endfunction 
  